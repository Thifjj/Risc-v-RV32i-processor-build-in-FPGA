library IEEE;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Rom_32bit is
	port(
		i_ADDR : in std_logic_vector(31 downto 0);
		o_INST : out std_logic_vector(31 downto 0)
	);
end entity Rom_32bit;

architecture arch of Rom_32bit is

	type T_ROM_ARRAY is array (0 to 255) of std_logic_vector(7 downto 0);
	constant ROM : T_ROM_ARRAY := (
	"00000001", "00000000", "00000100", "00010011",  -- addi s0, zero, 16
	"00000100", "00000000", "00000100", "10010011",  -- addi s9, zero, 64
	"00000000", "00010000", "00001001", "00010011",  -- addi s2, zero, 1
	"00000000", "00100000", "00001001", "10010011",  -- addi s3, zero, 2
	"00000000", "00110000", "00001010", "00010011",  -- addi a0, zero, 3
	"00000000", "01000000", "00001010", "10010011",  -- addi a1, zero, 4
	"00000000", "01010000", "00001011", "00010011",  -- addi a2, zero, 5
	"00000000", "01100000", "00001011", "10010011",  -- addi s7, zero, 6
	"00000000", "01110000", "00001100", "00010011",  -- addi a2, zero, 7
	"00000000", "10000000", "00001100", "10010011",  -- addi s9, zero, 8
	"00000000", "10010000", "00001101", "00010011",  -- addi a3, zero, 9
	"00000000", "10100000", "00001101", "10010011",  -- addi s11, zero, 10
	"00000000", "10110000", "00000011", "00010011",  -- addi t1, zero, 11
	"00000000", "11000000", "00000011", "10010011",  -- addi t2, zero, 12
	"00000000", "11010000", "00001110", "00010011",  -- addi a4, zero, 13
	"00000000", "11100000", "00001110", "10010011",  -- addi s9, zero, 14
	"00000000", "11110000", "00001111", "00010011",  -- addi a5, zero, 15
	"00000001", "00000000", "00001111", "10010011",  -- addi s3, zero, 16
	"00000000", "10010100", "00001001", "00110011",  -- add s2, s0, s1
	"00000001", "00111010", "00001010", "10110011",  -- add s5, s4, s3
	"00000001", "01101011", "10001100", "00110011",  -- add s8, s7, s6
	"00000001", "10101100", "10001101", "10110011",  -- add s11, s9, s8
	"01000000", "10010100", "10000100", "00110011",  -- sub s0, s1, s2
	"00000000", "00110000", "00000100", "10010011",  -- addi s9, zero, 3
	"00000000", "01000000", "00001001", "00010011",  -- addi s2, zero, 4
	"00000000", "01010000", "00001001", "10010011",  -- addi s3, zero, 5
	"00000000", "01100000", "00001010", "00010011",  -- addi a0, zero, 6
	"00000000", "01110000", "00001010", "10010011",  -- addi a1, zero, 7
	"00000000", "10000000", "00001011", "00010011",  -- addi a2, zero, 8
	"00000000", "10010000", "00001011", "10010011",  -- addi s7, zero, 9
	"00000000", "10100000", "00001100", "00010011",  -- addi a2, zero, 10
	"00000000", "10110000", "00001100", "10010011",  -- addi s9, zero, 11
	"00000000", "11000000", "00001101", "00010011",  -- addi a3, zero, 12
	"00000000", "00010000", "00000100", "10010011",  -- addi s9, zero, 1
	"00000000", "00100000", "00000100", "00010011",  -- addi s0, zero, 2
	"00000000", "00110000", "00000100", "10010011",  -- addi s9, zero, 3
		others => x"00"
	);
begin
o_INST <= ROM(to_integer(unsigned(i_ADDR))) &
ROM(to_integer(unsigned(i_ADDR))+1) &
ROM(to_integer(unsigned(i_ADDR))+2) &
ROM(to_integer(unsigned(i_ADDR))+3);
end arch;